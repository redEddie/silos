//Define level sensitive latch using UDP.
primitive latch(q, d, clock, clear);

//declarations
output q;
reg q; //q declared as reg
input d, clock, clear;

//sequential UDP initialization
//only one initial statement allowed
initial
    q = 0; 

//state table
table
  //d  clock  clear  : q  :  q+ ;
  
    ?    ?    1      :  ?  : 0  ;  //clear condition; 
                                   //q+ is the new output value
      
    1    1    0      :  ?  :  1 ; //latch q = data  = 1  
    0    1    0      :  ?  :  0 ; //latch q = data  = 0  

    ?    0    0      :  ?  :  - ; //retain original state if clock = 0
endtable

endprimitive
    
//This file must be simulated with the file
//"edge_dff.v". Please include both files in the
//project file.

module stimulus;

wire Q;
reg D, CLK, RESET;

always #5 CLK = ~CLK;

initial
begin
	$monitor($time, " Q=%b, D= %b, CLK=%b, RESET = %b",
			Q, D, CLK, RESET);
	RESET = 1'B1;
	CLK = 1'B0;
	#10 RESET = 1'B0;

	D = 1'b0;
	#110 D = 1'b0;
        #150 D = 1'b1;	
	#100 $stop;
end
 
//instantiate the d-flipflop
latch L(Q,  D, CLK, RESET);
 
endmodule
