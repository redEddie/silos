//This file cannot be simulated or compiled as a Verilog file.

The basic components of a module definition are:

1. Module, module name

2. port list

3. Parameters

4. Declarations of wires, regs and other variables

5. Instantiation of lower level modules

6. Data flow statements (assign)

7. always and initial blocks

8. tasks and functions

9. endmodule


All components except keyword module, module name and keyword endmodule
are optional.

