//This file does not really do anything.
//It only demonstrates the declaration of an integer.
module integer_example;

integer counter; // general purpose variable used as a counter.
initial
	counter = -1; // A negative one is stored in the counter

endmodule


